*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/RPLY_EX0_lpe.spi
#else
.include ../../../work/xsch/RPLY_EX0.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
IBP 0 IBPS_4U dc 4u
V0  IBNS_20U 0 dc 1

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VSS IBPS_4U IBNS_20U RPLY_EX0

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(VSS) v(IBPS_4U) v(IBNS_20U) i(V0)
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100p 2n 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
tran 10p 20n 1p
write
quit
#endif

.endc

.end
